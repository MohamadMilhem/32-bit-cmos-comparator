*** SPICE deck for cell PrefixAdderBased32bitComparatorNEW{lay} from library IC_PROJECT_FINAL_VERSION
*** Created on Sun Aug 18, 2024 20:37:09
*** Last revised on Thu Aug 22, 2024 18:28:41
*** Written on Thu Aug 22, 2024 18:49:45 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__Generate FROM CELL Generate{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__Generate g1 g2 gnd out p2 vdd
Mnmos@0 net@6 g1 gnd gnd NMOS L=0.044U W=0.352U AS=0.085P AD=0.025P PS=1.529U PD=0.836U
Mnmos@1 gnd g2 out gnd NMOS L=0.044U W=0.176U AS=0.055P AD=0.085P PS=1.085U PD=1.529U
Mnmos@2 out p2 net@6 gnd NMOS L=0.044U W=0.352U AS=0.025P AD=0.055P PS=0.836U PD=1.085U
Mpmos@0 net@0 p2 vdd vdd PMOS L=0.044U W=0.704U AS=0.12P AD=0.072P PS=1.892U PD=1.144U
Mpmos@1 vdd g1 net@0 vdd PMOS L=0.044U W=0.704U AS=0.072P AD=0.12P PS=1.144U PD=1.892U
Mpmos@2 net@0 g2 out vdd PMOS L=0.044U W=0.704U AS=0.055P AD=0.072P PS=1.085U PD=1.144U
.ENDS IC_PROJECT_FINAL_VERSION__Generate

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__inv FROM CELL inv{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__inv gnd in out vdd
Mnmos@0 gnd in out gnd NMOS L=0.044U W=0.176U AS=0.038P AD=0.078P PS=0.814U PD=1.826U
Mpmos@0 vdd in out vdd PMOS L=0.044U W=0.352U AS=0.038P AD=0.12P PS=0.814U PD=2.31U
.ENDS IC_PROJECT_FINAL_VERSION__inv

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__nand FROM CELL nand{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__nand A B gnd out vdd
Mnmos@0 net@20 B out gnd NMOS L=0.044U W=0.352U AS=0.043P AD=0.023P PS=0.711U PD=0.484U
Mnmos@1 gnd A net@20 gnd NMOS L=0.044U W=0.352U AS=0.023P AD=0.142P PS=0.484U PD=2.882U
Mpmos@0 out B vdd vdd PMOS L=0.044U W=0.352U AS=0.161P AD=0.043P PS=2.926U PD=0.711U
Mpmos@1 net@21 A out vdd PMOS L=0.044U W=0.352U AS=0.043P AD=0.058P PS=0.711U PD=1.034U
.ENDS IC_PROJECT_FINAL_VERSION__nand

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__PGNEW FROM CELL PGNEW{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__PGNEW g1 g2 Gi gnd p1 p2 Pi vdd
XGenerate@2 g1 g2 gnd net@192 p2 vdd IC_PROJECT_FINAL_VERSION__Generate
Xinv@6 gnd net@192 Gi vdd IC_PROJECT_FINAL_VERSION__inv
Xinv@7 gnd net@145 Pi vdd IC_PROJECT_FINAL_VERSION__inv
Xnand@3 p2 p1 gnd net@145 vdd IC_PROJECT_FINAL_VERSION__nand
.ENDS IC_PROJECT_FINAL_VERSION__PGNEW

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__xor FROM CELL xor{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__xor A B gnd out vdd
Xinv@0 gnd A out vdd IC_PROJECT_FINAL_VERSION__inv
Mnmos@0 gnd A A gnd NMOS L=0.044U W=0.176U AS=0.038P AD=0.025P PS=0.814U PD=0.638U
Mpmos@0 net@42 A A vdd PMOS L=0.044U W=0.352U AS=0.038P AD=0.031P PS=0.814U PD=0.528U
Mpmos@1 B B net@42 vdd PMOS L=0.044U W=0.352U AS=0.031P AD=0.05P PS=0.528U PD=0.99U
.ENDS IC_PROJECT_FINAL_VERSION__xor

*** SUBCIRCUIT IC_PROJECT_FINAL_VERSION__preifx_AdderNEW FROM CELL preifx_AdderNEW{lay}
.SUBCKT IC_PROJECT_FINAL_VERSION__preifx_AdderNEW Ai Bi GI gnd Pi vdd
Xinv@4 gnd Bi net@167 vdd IC_PROJECT_FINAL_VERSION__inv
Xinv@5 gnd net@185 GI vdd IC_PROJECT_FINAL_VERSION__inv
Xnand@3 net@167 Ai gnd net@185 vdd IC_PROJECT_FINAL_VERSION__nand
Xxor@3 Bi Ai gnd Pi vdd IC_PROJECT_FINAL_VERSION__xor
.ENDS IC_PROJECT_FINAL_VERSION__preifx_AdderNEW

*** TOP LEVEL CELL: PrefixAdderBased32bitComparatorNEW{lay}
XPGNEW@3 net@77 net@83 net@172 gnd ptest net@81 net@170 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@4 net@62 net@72 net@166 gnd net@64 net@69 net@159 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@5 net@166 net@172 net@2095 gnd net@159 net@170 net@2091 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@6 net@2431 net@2437 net@2501 gnd net@2429 net@2435 net@2499 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@7 net@2416 net@2426 net@2495 gnd net@2418 net@2423 net@2488 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@8 net@2495 net@2501 net@2519 gnd net@2488 net@2499 net@2516 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@9 net@2095 net@2519 net@3426 gnd net@2091 net@2516 net@3421 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@10 net@2586 net@2592 net@2656 gnd net@2584 net@2590 net@2654 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@11 net@2571 net@2581 net@2650 gnd net@2573 net@2578 net@2643 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@12 net@2650 net@2656 net@2674 gnd net@2643 net@2654 net@2671 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@13 net@2732 net@2738 net@2802 gnd net@2730 net@2736 net@2800 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@14 net@2717 net@2727 net@2796 gnd net@2719 net@2724 net@2789 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@15 net@2796 net@2802 net@2819 gnd net@2789 net@2800 net@2817 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@16 net@2674 net@2819 net@3435 gnd net@2671 net@2817 net@3438 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@31 net@3426 net@3435 net@4102 gnd net@3421 net@3438 net@4096 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@33 net@3509 net@3515 net@3579 gnd net@3507 net@3513 net@3577 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@34 net@3494 net@3504 net@3573 gnd net@3496 net@3501 net@3566 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@35 net@3573 net@3579 net@3597 gnd net@3566 net@3577 net@3594 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@36 net@3655 net@3661 net@3725 gnd net@3653 net@3659 net@3723 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@37 net@3640 net@3650 net@3719 gnd net@3642 net@3647 net@3712 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@38 net@3719 net@3725 net@3742 gnd net@3712 net@3723 net@3740 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@39 net@3597 net@3742 net@4052 gnd net@3594 net@3740 net@4047 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@40 net@3803 net@3809 net@3873 gnd net@3801 net@3807 net@3871 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@41 net@3788 net@3798 net@3867 gnd net@3790 net@3795 net@3860 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@42 net@3867 net@3873 net@3891 gnd net@3860 net@3871 net@3888 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@43 net@3949 net@3955 net@4019 gnd net@3947 net@3953 net@4017 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@44 net@3934 net@3944 net@4013 gnd net@3936 net@3941 net@4006 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@45 net@4013 net@4019 net@4036 gnd net@4006 net@4017 net@4034 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@46 net@3891 net@4036 net@4059 gnd net@3888 net@4034 net@4062 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@47 net@4052 net@4059 net@4079 gnd net@4047 net@4062 net@4077 vdd IC_PROJECT_FINAL_VERSION__PGNEW
XPGNEW@48 net@4102 net@4079 GT gnd net@4096 net@4077 EQ vdd IC_PROJECT_FINAL_VERSION__PGNEW
Xinv@0 gnd GT LT vdd IC_PROJECT_FINAL_VERSION__inv
Xpreifx_A@7 A0 B0 net@62 gnd net@64 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@8 A1 B1 net@72 gnd net@69 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@9 A2 B2 net@77 gnd ptest vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@10 A3 B3 net@83 gnd net@81 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@11 A4 B4 net@2416 gnd net@2418 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@12 A5 B5 net@2426 gnd net@2423 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@13 A6 B6 net@2431 gnd net@2429 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@14 A7 B7 net@2437 gnd net@2435 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@15 A8 B8 net@2571 gnd net@2573 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@16 A9 B9 net@2581 gnd net@2578 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@17 A10 B10 net@2586 gnd net@2584 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@18 A11 B11 net@2592 gnd net@2590 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@19 A12 B12 net@2717 gnd net@2719 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@20 A13 B13 net@2727 gnd net@2724 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@21 A14 B14 net@2732 gnd net@2730 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@22 A15 B15 net@2738 gnd net@2736 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@39 A16 B16 net@3494 gnd net@3496 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@40 A17 B17 net@3504 gnd net@3501 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@41 A18 B18 net@3509 gnd net@3507 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@42 A19 B19 net@3515 gnd net@3513 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@43 A20 B20 net@3640 gnd net@3642 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@44 A21 B21 net@3650 gnd net@3647 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@45 A22 B22 net@3655 gnd net@3653 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@46 A23 B23 net@3661 gnd net@3659 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@47 A24 B24 net@3788 gnd net@3790 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@48 A25 B25 net@3798 gnd net@3795 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@49 A26 B26 net@3803 gnd net@3801 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@50 A27 B27 net@3809 gnd net@3807 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@51 A28 B28 net@3934 gnd net@3936 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@52 A29 B29 net@3944 gnd net@3941 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@53 A30 B30 net@3949 gnd net@3947 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW
Xpreifx_A@54 A31 B31 net@3955 gnd net@3953 vdd IC_PROJECT_FINAL_VERSION__preifx_AdderNEW

* Spice Code nodes in cell cell 'PrefixAdderBased32bitComparatorNEW{lay}'
Vdd vdd 0 DC 1.9
V_A0 A0 0 pwl 0n 0 22n 0 24n 1.9 46n 1.9 48n 0
V_A1 A1 0 DC 0
V_A2 A2 0 DC 0
V_A3 A3 0 DC 0
V_A4 A4 0 DC 0
V_A5 A5 0 DC 0
V_A6 A6 0 DC 0
V_A7 A7 0 DC 0
V_A8 A8 0 DC 0
V_A9 A9 0 DC 0
V_A10 A10 0 DC 0
V_A11 A11 0 DC 0
V_A12 A12 0 DC 0
V_A13 A13 0 DC 0
V_A14 A14 0 DC 1.9
V_A15 A15 0 DC 0
V_A16 A16 0 DC 0
V_A17 A17 0 DC 0
V_A18 A18 0 DC 0
V_A19 A19 0 DC 0
V_A20 A20 0 DC 0
V_A21 A21 0 DC 0
V_A22 A22 0 DC 0
V_A23 A23 0 DC 0
V_A24 A24 0 DC 0
V_A25 A25 0 DC 0
V_A26 A26 0 DC 0
V_A27 A27 0 DC 0
V_A28 A28 0 DC 0
V_A29 A29 0 DC 1.9
V_A30 A30 0 DC 1.9
V_A31 A31 0 DC 0
V_B0 B0 0 pwl 0n 0 10n 0 12n 1.9 22n 1.9 24n 0 34n 0 36n 1.9 46n 1.9 48n 0
V_B1 B1 0 DC 0
V_B2 B2 0 DC 0
V_B3 B3 0 DC 0
V_B4 B4 0 DC 0
V_B5 B5 0 DC 0
V_B6 B6 0 DC 0
V_B7 B7 0 DC 0
V_B8 B8 0 DC 0
V_B9 B9 0 DC 0
V_B10 B10 0 DC 0
V_B11 B11 0 DC 0
V_B12 B12 0 DC 0
V_B13 B13 0 DC 0
V_B14 B14 0 DC 1.9
V_B15 B15 0 DC 0
V_B16 B16 0 DC 0
V_B17 B17 0 DC 0
V_B18 B18 0 DC 0
V_B19 B19 0 DC 0
V_B20 B20 0 DC 0
V_B21 B21 0 DC 0
V_B22 B22 0 DC 0
V_B23 B23 0 DC 0
V_B24 B24 0 DC 0
V_B25 B25 0 DC 0
V_B26 B26 0 DC 0
V_B27 B27 0 DC 0
V_B28 B28 0 DC 0
V_B29 B29 0 DC 1.9
V_B30 B30 0 DC 1.9
V_B31 B31 0 DC 0
Cload_case11 GT 0 250fF
Cload_case12 LT 0 250fF
Cload_case13 EQ 0 250fF
.tran 0 60ns
.INCLUDE C:\22nm.txt
.END
